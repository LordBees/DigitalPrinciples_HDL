--dffasync